`ifndef TURFIO_DEBUG_VH
`define TURFIO_DEBUG_VH

`define TURF_INTERFACE_DEBUG "FALSE"
`define TURF_CIN_PARALLEL_SYNC_DEBUG "TRUE"

`endif
